library ieee;
   use ieee.std_logic_1164.all;


package wbfbd is

type t_slv_vector is array (natural range <>) of std_logic_vector;

-- Packages constants
{{.PkgsConsts}}
end package;
