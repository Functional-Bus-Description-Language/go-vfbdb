library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;

library ltypes;
   use ltypes.types.all;


package wb3 is

-- Packages constants
{{.PkgsConsts}}

end package;
