library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;

library types;
   use types.types.all;


package wbfbd is

-- Packages constants
{{.PkgsConsts}}

end package;
